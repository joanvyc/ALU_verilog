module nbit_shift #(parameter bits=8) (
	input [bits-1:0] A,
	input [$clog2(bits):0] B,
	output [bits-1:0] X);

	
endmodule
			